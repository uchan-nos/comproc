`define ADDR_WIDTH 12
