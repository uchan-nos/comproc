`define ADDR_WIDTH 10
